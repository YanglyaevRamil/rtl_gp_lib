//***************  ****************************


//**************************************************************